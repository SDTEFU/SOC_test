// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : fetch_mem
// Git hash  : c4ec9e181b11aa1052ddd4f4a0813de50e3648a5

`timescale 1ns/1ps

module fetch_mem (
  input               io_ex_en,
  input               io_ex_w_en,
  input      [31:0]   io_ex_mem_addr,
  input               io_SSE_belong,
  input               io_SSE_done
);



endmodule
