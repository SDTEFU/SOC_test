// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : template_module
// Git hash  : 232a2cb27d43b74a1342826f9bbd0f790b781192

`timescale 1ns/1ps

module template_module (
);



endmodule
