// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : temp
// Git hash  : d1c9adfb9a7aab45a29ba6b84e3bea900a8c7bee

`timescale 1ns/1ps

module temp (
);



endmodule
