// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : temp
// Git hash  : dc2fba5c92e024ce30402f160bd755ad38650a3b

`timescale 1ns/1ps

module temp (
);



endmodule
