// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : temp
// Git hash  : c4ec9e181b11aa1052ddd4f4a0813de50e3648a5

`timescale 1ns/1ps

module temp (
);



endmodule
