// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : IFetch
// Git hash  : 8c6c7cf9176f84e124a944713de8a584b5d63265

`timescale 1ns/1ps

module IFetch (
);



endmodule
