// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : temp
// Git hash  : 4fb0decdf9108ab8284140c032b988fb222abb89

`timescale 1ns/1ps

module temp (
);



endmodule
