// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : IFetch
// Git hash  : 42245be0c103b6f7a97635b2c19f9bae38093db0

`timescale 1ns/1ps

module IFetch (
);



endmodule
