// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : IFetch
// Git hash  : 54169215138359a268c1d14a644c4d66f6ca19d3

`timescale 1ns/1ps

module IFetch (
);



endmodule
